LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
USE ieee.std_logic_unsigned.ALL;
use IEEE.std_logic_arith.all;

ENTITY SENSOR_CONTROL IS
	PORT(	ECHO, CLOCK	:	IN	STD_LOGIC;
			TRIG			:	OUT STD_LOGIC; -- RECEIVE FROM ECHO PIN
			OUT1, OUT2	:	OUT STD_LOGIC; -- CONTROL
			EN				:	IN STD_LOGIC -- ENABLE WHICH CONTROL
			);
END ENTITY;

ARCHITECTURE CONTROL OF SENSOR_CONTROL IS
BEGIN

PROCESS(CLOCK)
VARIABLE COUNT1, COUNT2	: INTEGER	:= 0; -- COUNT CLOCK CYCLE
VARIABLE ECHO_COUNT		: INTEGER	:= 0; -- CALCULATE DISTANCE
VARIABLE MASK				: STD_LOGIC	:= '1';	
BEGIN
	IF(EN = '1') THEN
		IF(RISING_EDGE(CLOCK)) THEN
			--INPUTTING SIGNAL
			IF (COUNT1 = 0) THEN -- START GIVING OUT SIGNAL HIGH
				TRIG <= '1';
			ELSIF(COUNT1 = 500) THEN -- COUNT UP TO 10 US
				TRIG <= '0'; -- DONE OUTPUTTING SIGNAL
				MASK	:= '1';
			ELSIF(COUNT1 = 5000000) THEN -- COUNT UP TO 100 MS
				TRIG <= '1';
				COUNT1 := 0; -- RESET COUNTER
			END IF;
			COUNT1 := COUNT1 + 1; -- INCREASE THE COUNTER
			
			--DETECT ECHO
			IF(ECHO = '1') THEN
				COUNT2 := COUNT2 + 1;
			ELSIF(ECHO = '0' AND MASK = '1') THEN
				ECHO_COUNT	:= COUNT2; 
				COUNT2	 	:= 0;	
				MASK			:= '0';
			END IF;
			
			--MAP THE GAME
			--USE THE FORMULA 1 US = 58*1 CM
			IF(ECHO_COUNT <= 58000) THEN -- IF THE DISTANCE LESS THAN 5 CM
				OUT1	<= '1'; -- MOVE POSITIVE DIRECTION
				OUT2	<= '0';
			ELSIF(ECHO_COUNT	> 58000) THEN-- IF THE DISTANCE BETWEEN 10CM AND 15 CM
				OUT1	<= '0';	-- MOVE NEGATIVE DIRECTION
				OUT2	<=	'1';
			ELSE
				OUT1	<= '0'; --STOP
				OUT2	<= '0';
			END IF;
		END IF;
	ELSE
		TRIG <= '0';
		OUT1 <= '0';
		OUT2 <= '0';
		COUNT1 := 0;
		COUNT2 := 0;
	END IF;
END PROCESS;
END CONTROL;